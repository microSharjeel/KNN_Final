`timescale 1ns/1ps
`include "iob_lib.vh"
`include "interconnect.vh"
`include "iob_knn.vh"

module iob_knn
  #(
    parameter ADDR_W = `KNN_ADDR_W, 
    parameter DATA_W = 32, 
    parameter WDATA_W = `KNN_WDATA_W 
    )
	(
	//CPU native interface	
	//cpu generic slave interface copied from
	`include "cpu_nat_s_if.v"
	//clk rst generic interface copied from
	`include "gen_if.v"
	);
	`include "KNN_Header.vh"
 	`include "KNNsw_reg.v"
	`include "KNNsw_reg_gen.v"

	`SIGNAL_OUT(KNN_VALID_OUT_TOP,1)
	`SIGNAL_OUT(KN1_OUT_TOP,`WDATA_W)
	`SIGNAL_OUT(KN2_OUT_TOP,`WDATA_W)
	`SIGNAL_OUT(KN3_OUT_TOP,`WDATA_W)
	`SIGNAL_OUT(KN4_OUT_TOP,`WDATA_W)
	`SIGNAL_OUT(KN5_OUT_TOP,`WDATA_W)
	`SIGNAL_OUT(KN6_OUT_TOP,`WDATA_W)
	
	`SIGNAL_OUT(IN1_OUT_TOP,`K_NUM_DATA_PTS_BIT)
	`SIGNAL_OUT(IN2_OUT_TOP,`K_NUM_DATA_PTS_BIT)
	`SIGNAL_OUT(IN3_OUT_TOP,`K_NUM_DATA_PTS_BIT)
	`SIGNAL_OUT(IN4_OUT_TOP,`K_NUM_DATA_PTS_BIT)
	`SIGNAL_OUT(IN5_OUT_TOP,`K_NUM_DATA_PTS_BIT)
	`SIGNAL_OUT(IN6_OUT_TOP,`K_NUM_DATA_PTS_BIT)
	
	wire rst_comb;
	assign rst_comb = rst | KNN_RESET;
	/* 
	knn_core  knn_core_top
	 (
	  .KNN_START_CORE    (KNN_START),
	  .KNN_DATA_PT_CORE1  (KNN_DATA_PT1), 
	  .KNN_DATA_PT_CORE2  (KNN_DATA_PT2), 
	  .KNN_DATA_PT_CORE3  (KNN_DATA_PT3), 
	  .KNN_DATA_PT_CORE4  (KNN_DATA_PT4), 
  	  .KNN_DATA_PT_CORE5  (KNN_DATA_PT5), 
	  .KNN_DATA_PT_CORE6  (KNN_DATA_PT6), 
	  .KNN_DATA_PT_CORE7  (KNN_DATA_PT7), 
	  .KNN_DATA_PT_CORE8  (KNN_DATA_PT8), 
	  .KNN_TEST_PT_CORE  (KNN_TEST_PT),
	  .KNN_VALID_CORE    (KNN_VALID_IN),
	  .KNN_SAMPLE_CORE   (KNN_SAMPLE),
	  .KNN_VALID_OUT_CORE(KNN_VALID_OUT_TOP),
	 
	  .KN1_OUT_CORE(KN1_OUT_TOP),
	  .KN2_OUT_CORE(KN2_OUT_TOP),
	  .KN3_OUT_CORE(KN3_OUT_TOP),
	  .KN4_OUT_CORE(KN4_OUT_TOP),
	  .KN5_OUT_CORE(KN5_OUT_TOP),
	  .KN6_OUT_CORE(KN6_OUT_TOP),

	  .IN1_OUT_CORE(IN1_OUT_TOP),
	  .IN2_OUT_CORE(IN2_OUT_TOP),
	  .IN3_OUT_CORE(IN3_OUT_TOP),
	  .IN4_OUT_CORE(IN4_OUT_TOP),
	  .IN5_OUT_CORE(IN5_OUT_TOP),
	  .IN6_OUT_CORE(IN6_OUT_TOP),

	  .CLK_CORE(clk),
	  .RST_CORE(rst_comb)

	 );
*/

//////////////////////////////////////
knn_core knn_core_top

(
  .KNN_START_CORE    (KNN_START),

  .KNN_DATA_PT_CORE0  (KNN_DATA_PT0), 
  .KNN_DATA_PT_CORE1  (KNN_DATA_PT1), 
  .KNN_DATA_PT_CORE2  (KNN_DATA_PT2), 
  .KNN_DATA_PT_CORE3  (KNN_DATA_PT3), 
  .KNN_DATA_PT_CORE4  (KNN_DATA_PT4), 
  .KNN_DATA_PT_CORE5  (KNN_DATA_PT5), 
  .KNN_DATA_PT_CORE6  (KNN_DATA_PT6), 
  .KNN_DATA_PT_CORE7  (KNN_DATA_PT7), 

  .KNN_DATA_PT_CORE8  (KNN_DATA_PT8), 
  .KNN_DATA_PT_CORE9  (KNN_DATA_PT9), 
  .KNN_DATA_PT_CORE10  (KNN_DATA_PT10), 
  .KNN_DATA_PT_CORE11  (KNN_DATA_PT11), 
  .KNN_DATA_PT_CORE12  (KNN_DATA_PT12), 
  .KNN_DATA_PT_CORE13  (KNN_DATA_PT13), 
  .KNN_DATA_PT_CORE14  (KNN_DATA_PT14), 
  .KNN_DATA_PT_CORE15  (KNN_DATA_PT15), 

  .KNN_DATA_PT_CORE16  (KNN_DATA_PT16), 
  .KNN_DATA_PT_CORE17  (KNN_DATA_PT17), 
  .KNN_DATA_PT_CORE18  (KNN_DATA_PT18), 
  .KNN_DATA_PT_CORE19  (KNN_DATA_PT19), 
  .KNN_DATA_PT_CORE20  (KNN_DATA_PT20), 
  .KNN_DATA_PT_CORE21  (KNN_DATA_PT21), 
  .KNN_DATA_PT_CORE22  (KNN_DATA_PT22), 
  .KNN_DATA_PT_CORE23  (KNN_DATA_PT23),
  
  
  .KNN_DATA_PT_CORE24  (KNN_DATA_PT24), 
  .KNN_DATA_PT_CORE25  (KNN_DATA_PT25), 
  .KNN_DATA_PT_CORE26  (KNN_DATA_PT26), 
  .KNN_DATA_PT_CORE27  (KNN_DATA_PT27), 
  .KNN_DATA_PT_CORE28  (KNN_DATA_PT28), 
  .KNN_DATA_PT_CORE29  (KNN_DATA_PT29), 
  .KNN_DATA_PT_CORE30  (KNN_DATA_PT30), 
  .KNN_DATA_PT_CORE31  (KNN_DATA_PT31),
  
  
  .KNN_DATA_PT_CORE32  (KNN_DATA_PT32), 
  .KNN_DATA_PT_CORE33  (KNN_DATA_PT33), 
  .KNN_DATA_PT_CORE34  (KNN_DATA_PT34), 
  .KNN_DATA_PT_CORE35  (KNN_DATA_PT35), 
  .KNN_DATA_PT_CORE36  (KNN_DATA_PT36), 
  .KNN_DATA_PT_CORE37  (KNN_DATA_PT37), 
  .KNN_DATA_PT_CORE38  (KNN_DATA_PT38), 
  .KNN_DATA_PT_CORE39  (KNN_DATA_PT39),
  
  .KNN_DATA_PT_CORE40  (KNN_DATA_PT40), 
  .KNN_DATA_PT_CORE41  (KNN_DATA_PT41), 
  .KNN_DATA_PT_CORE42  (KNN_DATA_PT42), 
  .KNN_DATA_PT_CORE43  (KNN_DATA_PT43), 
  .KNN_DATA_PT_CORE44  (KNN_DATA_PT44), 
  .KNN_DATA_PT_CORE45  (KNN_DATA_PT45), 
  .KNN_DATA_PT_CORE46  (KNN_DATA_PT46), 
  .KNN_DATA_PT_CORE47  (KNN_DATA_PT47),

  .KNN_DATA_PT_CORE48  (KNN_DATA_PT48),
  .KNN_DATA_PT_CORE49  (KNN_DATA_PT49), 
  .KNN_DATA_PT_CORE50  (KNN_DATA_PT50), 
  .KNN_DATA_PT_CORE51  (KNN_DATA_PT51), 
  .KNN_DATA_PT_CORE52  (KNN_DATA_PT52), 
  .KNN_DATA_PT_CORE53  (KNN_DATA_PT53), 
  .KNN_DATA_PT_CORE54  (KNN_DATA_PT54), 
  .KNN_DATA_PT_CORE55  (KNN_DATA_PT55), 

  .KNN_DATA_PT_CORE56  (KNN_DATA_PT56),
  
  .KNN_DATA_PT_CORE57  (KNN_DATA_PT57), 
  .KNN_DATA_PT_CORE58  (KNN_DATA_PT58), 
  .KNN_DATA_PT_CORE59  (KNN_DATA_PT59), 
  .KNN_DATA_PT_CORE60  (KNN_DATA_PT60), 
  .KNN_DATA_PT_CORE61  (KNN_DATA_PT61), 
  .KNN_DATA_PT_CORE62  (KNN_DATA_PT62), 
  .KNN_DATA_PT_CORE63  (KNN_DATA_PT63), 
  .KNN_DATA_PT_CORE64  (KNN_DATA_PT64),
  
  .KNN_DATA_PT_CORE65  (KNN_DATA_PT65), 
  .KNN_DATA_PT_CORE66  (KNN_DATA_PT66), 
  .KNN_DATA_PT_CORE67  (KNN_DATA_PT67), 
  .KNN_DATA_PT_CORE68  (KNN_DATA_PT68), 
  .KNN_DATA_PT_CORE69  (KNN_DATA_PT69), 
  .KNN_DATA_PT_CORE70  (KNN_DATA_PT70), 
  .KNN_DATA_PT_CORE71  (KNN_DATA_PT71), 
  .KNN_DATA_PT_CORE72  (KNN_DATA_PT72),
  
  .KNN_DATA_PT_CORE73  (KNN_DATA_PT73), 
  .KNN_DATA_PT_CORE74  (KNN_DATA_PT74), 
  .KNN_DATA_PT_CORE75  (KNN_DATA_PT75), 
  .KNN_DATA_PT_CORE76  (KNN_DATA_PT76), 
  .KNN_DATA_PT_CORE77  (KNN_DATA_PT77), 
  .KNN_DATA_PT_CORE78  (KNN_DATA_PT78), 
  .KNN_DATA_PT_CORE79  (KNN_DATA_PT79), 
  .KNN_DATA_PT_CORE80  (KNN_DATA_PT80),
  
  .KNN_DATA_PT_CORE81  (KNN_DATA_PT81), 
  .KNN_DATA_PT_CORE82  (KNN_DATA_PT82), 
  .KNN_DATA_PT_CORE83  (KNN_DATA_PT83), 
  .KNN_DATA_PT_CORE84  (KNN_DATA_PT84), 
  .KNN_DATA_PT_CORE85  (KNN_DATA_PT85), 
  .KNN_DATA_PT_CORE86  (KNN_DATA_PT86), 
  .KNN_DATA_PT_CORE87  (KNN_DATA_PT87), 
  .KNN_DATA_PT_CORE88  (KNN_DATA_PT88),
  
  .KNN_DATA_PT_CORE89  (KNN_DATA_PT89), 
  .KNN_DATA_PT_CORE90  (KNN_DATA_PT90), 
  .KNN_DATA_PT_CORE91  (KNN_DATA_PT91), 
  .KNN_DATA_PT_CORE92  (KNN_DATA_PT92), 
  .KNN_DATA_PT_CORE93  (KNN_DATA_PT93), 
  .KNN_DATA_PT_CORE94  (KNN_DATA_PT94), 
  .KNN_DATA_PT_CORE95  (KNN_DATA_PT95), 
  .KNN_DATA_PT_CORE96  (KNN_DATA_PT96),
  
  
  .KNN_DATA_PT_CORE97  (KNN_DATA_PT97), 
  .KNN_DATA_PT_CORE98  (KNN_DATA_PT98), 
  .KNN_DATA_PT_CORE99  (KNN_DATA_PT99), 
  .KNN_DATA_PT_CORE100  (KNN_DATA_PT100), 
  .KNN_DATA_PT_CORE101  (KNN_DATA_PT101), 
  .KNN_DATA_PT_CORE102  (KNN_DATA_PT102), 
  .KNN_DATA_PT_CORE103  (KNN_DATA_PT103), 
  .KNN_DATA_PT_CORE104  (KNN_DATA_PT104),
  
  .KNN_DATA_PT_CORE105  (KNN_DATA_PT105), 
  .KNN_DATA_PT_CORE106  (KNN_DATA_PT106), 
  .KNN_DATA_PT_CORE107  (KNN_DATA_PT107), 
  .KNN_DATA_PT_CORE108  (KNN_DATA_PT108), 
  .KNN_DATA_PT_CORE109  (KNN_DATA_PT109), 
  .KNN_DATA_PT_CORE110  (KNN_DATA_PT110), 
  .KNN_DATA_PT_CORE111  (KNN_DATA_PT111), 
  .KNN_DATA_PT_CORE112  (KNN_DATA_PT112),
  
  .KNN_DATA_PT_CORE113  (KNN_DATA_PT113), 
  .KNN_DATA_PT_CORE114  (KNN_DATA_PT114), 
  .KNN_DATA_PT_CORE115  (KNN_DATA_PT115), 
  .KNN_DATA_PT_CORE116  (KNN_DATA_PT116), 
  .KNN_DATA_PT_CORE117  (KNN_DATA_PT117), 
  .KNN_DATA_PT_CORE118  (KNN_DATA_PT118), 
  .KNN_DATA_PT_CORE119  (KNN_DATA_PT119), 
  .KNN_DATA_PT_CORE120  (KNN_DATA_PT120),
  
  
  .KNN_DATA_PT_CORE121  (KNN_DATA_PT121), 
  .KNN_DATA_PT_CORE122  (KNN_DATA_PT122), 
  .KNN_DATA_PT_CORE123  (KNN_DATA_PT123), 
  .KNN_DATA_PT_CORE124  (KNN_DATA_PT124), 
  .KNN_DATA_PT_CORE125  (KNN_DATA_PT125), 
  .KNN_DATA_PT_CORE126  (KNN_DATA_PT126), 
  .KNN_DATA_PT_CORE127  (KNN_DATA_PT127), 
  
  
  .KNN_TEST_PT_CORE  (KNN_TEST_PT),
  .KNN_VALID_CORE    (KNN_VALID_IN),
  .KNN_SAMPLE_CORE   (KNN_SAMPLE),
  .KNN_VALID_OUT_CORE(KNN_VALID_OUT_TOP),
	 
  .KN1_OUT_CORE(KN1_OUT_TOP),
  .KN2_OUT_CORE(KN2_OUT_TOP),
  .KN3_OUT_CORE(KN3_OUT_TOP),
  .KN4_OUT_CORE(KN4_OUT_TOP),
  .KN5_OUT_CORE(KN5_OUT_TOP),
  .KN6_OUT_CORE(KN6_OUT_TOP),

  .IN1_OUT_CORE(IN1_OUT_TOP),
  .IN2_OUT_CORE(IN2_OUT_TOP),
  .IN3_OUT_CORE(IN3_OUT_TOP),
  .IN4_OUT_CORE(IN4_OUT_TOP),
  .IN5_OUT_CORE(IN5_OUT_TOP),
  .IN6_OUT_CORE(IN6_OUT_TOP),

  .CLK_CORE(clk),
  .RST_CORE(rst_comb)


);

/////////////////////////////////////////
	assign KNN_VALID_OUT = KNN_VALID_OUT_TOP;
	assign KNN_KN1 = KN1_OUT_TOP;
	assign KNN_KN2 = KN2_OUT_TOP;
	assign KNN_KN3 = KN3_OUT_TOP;
	assign KNN_KN4 = KN4_OUT_TOP;
	assign KNN_KN5 = KN5_OUT_TOP;
	assign KNN_KN6 = KN6_OUT_TOP;
	
	assign KNN_IN1 = IN1_OUT_TOP;
	assign KNN_IN2 = IN2_OUT_TOP;
	assign KNN_IN3 = IN3_OUT_TOP;
	assign KNN_IN4 = IN4_OUT_TOP;
	assign KNN_IN5 = IN5_OUT_TOP;
	assign KNN_IN6 = IN6_OUT_TOP;

		
endmodule
