`timescale 1ns/1ps
`include "KNN_Header.vh"
`include "iob_lib.vh"
 module knn_core
(
  `INPUT(KNN_START_CORE,1),
  `INPUT(KNN_DATA_PT_CORE0,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE1,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE2,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE3,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE4,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE5,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE6,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE7,`WDATA_W),
  
  `INPUT(KNN_DATA_PT_CORE8,`WDATA_W),  
  `INPUT(KNN_DATA_PT_CORE9,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE10,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE11,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE12,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE13,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE14,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE15,`WDATA_W),

  
  `INPUT(KNN_DATA_PT_CORE16,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE17,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE18,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE19,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE20,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE21,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE22,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE23,`WDATA_W),
  
  `INPUT(KNN_DATA_PT_CORE24,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE25,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE26,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE27,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE28,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE29,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE30,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE31,`WDATA_W),
  
  `INPUT(KNN_DATA_PT_CORE32,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE33,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE34,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE35,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE36,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE37,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE38,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE39,`WDATA_W),
  
  `INPUT(KNN_DATA_PT_CORE40,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE41,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE42,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE43,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE44,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE45,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE46,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE47,`WDATA_W),
  
  
  `INPUT(KNN_DATA_PT_CORE48,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE49,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE50,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE51,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE52,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE53,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE54,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE55,`WDATA_W),
  
  `INPUT(KNN_DATA_PT_CORE56,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE57,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE58,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE59,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE60,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE61,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE62,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE63,`WDATA_W),
  
  `INPUT(KNN_DATA_PT_CORE64,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE65,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE66,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE67,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE68,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE69,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE70,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE71,`WDATA_W),
  
  `INPUT(KNN_DATA_PT_CORE72,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE73,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE74,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE75,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE76,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE77,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE78,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE79,`WDATA_W),
  
  `INPUT(KNN_DATA_PT_CORE80,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE81,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE82,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE83,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE84,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE85,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE86,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE87,`WDATA_W),
  
  `INPUT(KNN_DATA_PT_CORE88,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE89,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE90,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE91,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE92,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE93,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE94,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE95,`WDATA_W),
  
  
  `INPUT(KNN_DATA_PT_CORE96,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE97,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE98,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE99,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE100,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE101,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE102,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE103,`WDATA_W),
  
  `INPUT(KNN_DATA_PT_CORE104,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE105,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE106,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE107,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE108,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE109,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE110,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE111,`WDATA_W),
  
  `INPUT(KNN_DATA_PT_CORE112,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE113,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE114,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE115,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE116,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE117,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE118,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE119,`WDATA_W),
  
  
  `INPUT(KNN_DATA_PT_CORE120,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE121,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE122,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE123,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE124,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE125,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE126,`WDATA_W),
  `INPUT(KNN_DATA_PT_CORE127,`WDATA_W),
  
  
  `INPUT(KNN_TEST_PT_CORE,`WDATA_W),
  `INPUT(KNN_VALID_CORE,1),
  `INPUT(KNN_SAMPLE_CORE,1),
  `OUTPUT(KNN_VALID_OUT_CORE,1),
 
  `OUTPUT(KN1_OUT_CORE,`WDATA_W),
  `OUTPUT(KN2_OUT_CORE,`WDATA_W),
  `OUTPUT(KN3_OUT_CORE,`WDATA_W),
  `OUTPUT(KN4_OUT_CORE,`WDATA_W),
  `OUTPUT(KN5_OUT_CORE,`WDATA_W),
  `OUTPUT(KN6_OUT_CORE,`WDATA_W),

  `OUTPUT(IN1_OUT_CORE,`K_NUM_DATA_PTS_BIT),
  `OUTPUT(IN2_OUT_CORE,`K_NUM_DATA_PTS_BIT),
  `OUTPUT(IN3_OUT_CORE,`K_NUM_DATA_PTS_BIT),
  `OUTPUT(IN4_OUT_CORE,`K_NUM_DATA_PTS_BIT),
  `OUTPUT(IN5_OUT_CORE,`K_NUM_DATA_PTS_BIT),
  `OUTPUT(IN6_OUT_CORE,`K_NUM_DATA_PTS_BIT),

  `INPUT(CLK_CORE, 1),
  `INPUT(RST_CORE, 1)

);

`SIGNAL_OUT(KNN_TST_CORE,`WDATA_W)
`SIGNAL_OUT(KNN_DAT_CORE,`WDATA_W)
`SIGNAL_OUT(KNN_ST_CORE,1)
/*
knn_fsm  knn_fsm_inst
(
	//to and from datapath
	.KNN_TEST_PT_O    (KNN_TST_CORE),
	.KNN_DATA_PT_O    (KNN_DAT_CORE),
	.KNN_START_O      (KNN_ST_CORE),
	//to and from KNN top level and KNN core 
	.KNN_START_FSM    (KNN_START_CORE),
	.KNN_DATA_PT_FSM1  (KNN_DATA_PT_CORE1),
	.KNN_DATA_PT_FSM2  (KNN_DATA_PT_CORE2),
	.KNN_DATA_PT_FSM3  (KNN_DATA_PT_CORE3),
	.KNN_DATA_PT_FSM4  (KNN_DATA_PT_CORE4),
	.KNN_DATA_PT_FSM5  (KNN_DATA_PT_CORE5),
	.KNN_DATA_PT_FSM6  (KNN_DATA_PT_CORE6),
	.KNN_DATA_PT_FSM7  (KNN_DATA_PT_CORE7),
	.KNN_DATA_PT_FSM8  (KNN_DATA_PT_CORE8),
	.KNN_TEST_PT_FSM  (KNN_TEST_PT_CORE),
	.KNN_VALID_IN_FSM (KNN_VALID_CORE),
	.KNN_VALID_O      (KNN_VALID_OUT_CORE),
	.clk(CLK_CORE),
	.rst(RST_CORE)
);
*/
knn_fsm  knn_fsm_inst

(
	//to and from datapath
	.KNN_TEST_PT_O    (KNN_TST_CORE),
	.KNN_DATA_PT_O    (KNN_DAT_CORE),
	.KNN_START_O      (KNN_ST_CORE),
	//to and from KNN top level and KNN core 
	.KNN_START_FSM    (KNN_START_CORE),
	.KNN_DATA_PT_FSM0  (KNN_DATA_PT_CORE0),
	.KNN_DATA_PT_FSM1  (KNN_DATA_PT_CORE1),
	.KNN_DATA_PT_FSM2  (KNN_DATA_PT_CORE2),
	.KNN_DATA_PT_FSM3  (KNN_DATA_PT_CORE3),
	.KNN_DATA_PT_FSM4  (KNN_DATA_PT_CORE4),
	.KNN_DATA_PT_FSM5  (KNN_DATA_PT_CORE5),
	.KNN_DATA_PT_FSM6  (KNN_DATA_PT_CORE6),
	.KNN_DATA_PT_FSM7  (KNN_DATA_PT_CORE7),
	
	.KNN_DATA_PT_FSM8  (KNN_DATA_PT_CORE8),
	.KNN_DATA_PT_FSM9  (KNN_DATA_PT_CORE9),
	.KNN_DATA_PT_FSM10  (KNN_DATA_PT_CORE10),
	.KNN_DATA_PT_FSM11  (KNN_DATA_PT_CORE11),
	.KNN_DATA_PT_FSM12  (KNN_DATA_PT_CORE12),
	.KNN_DATA_PT_FSM13  (KNN_DATA_PT_CORE13),
	.KNN_DATA_PT_FSM14  (KNN_DATA_PT_CORE14),
	.KNN_DATA_PT_FSM15  (KNN_DATA_PT_CORE15),
	
	
	.KNN_DATA_PT_FSM16  (KNN_DATA_PT_CORE16),
	.KNN_DATA_PT_FSM17  (KNN_DATA_PT_CORE17),
	.KNN_DATA_PT_FSM18  (KNN_DATA_PT_CORE18),
	.KNN_DATA_PT_FSM19  (KNN_DATA_PT_CORE19),
	.KNN_DATA_PT_FSM20  (KNN_DATA_PT_CORE20),
	.KNN_DATA_PT_FSM21  (KNN_DATA_PT_CORE21),
	.KNN_DATA_PT_FSM22  (KNN_DATA_PT_CORE22),
	.KNN_DATA_PT_FSM23  (KNN_DATA_PT_CORE23),
	
		
	.KNN_DATA_PT_FSM24  (KNN_DATA_PT_CORE24),
	.KNN_DATA_PT_FSM25  (KNN_DATA_PT_CORE25),
	.KNN_DATA_PT_FSM26  (KNN_DATA_PT_CORE26),
	.KNN_DATA_PT_FSM27  (KNN_DATA_PT_CORE27),
	.KNN_DATA_PT_FSM28  (KNN_DATA_PT_CORE28),
	.KNN_DATA_PT_FSM29  (KNN_DATA_PT_CORE29),
	.KNN_DATA_PT_FSM30  (KNN_DATA_PT_CORE30),
	.KNN_DATA_PT_FSM31  (KNN_DATA_PT_CORE31),
	
		
	.KNN_DATA_PT_FSM32  (KNN_DATA_PT_CORE32),
	.KNN_DATA_PT_FSM33  (KNN_DATA_PT_CORE33),
	.KNN_DATA_PT_FSM34  (KNN_DATA_PT_CORE34),
	.KNN_DATA_PT_FSM35  (KNN_DATA_PT_CORE35),
	.KNN_DATA_PT_FSM36  (KNN_DATA_PT_CORE36),
	.KNN_DATA_PT_FSM37  (KNN_DATA_PT_CORE37),
	.KNN_DATA_PT_FSM38  (KNN_DATA_PT_CORE38),
	.KNN_DATA_PT_FSM39  (KNN_DATA_PT_CORE39),
	
	.KNN_DATA_PT_FSM40  (KNN_DATA_PT_CORE40),
	.KNN_DATA_PT_FSM41  (KNN_DATA_PT_CORE41),
	.KNN_DATA_PT_FSM42  (KNN_DATA_PT_CORE42),
	.KNN_DATA_PT_FSM43  (KNN_DATA_PT_CORE43),
	.KNN_DATA_PT_FSM44  (KNN_DATA_PT_CORE44),
	.KNN_DATA_PT_FSM45  (KNN_DATA_PT_CORE45),
	.KNN_DATA_PT_FSM46  (KNN_DATA_PT_CORE46),
	.KNN_DATA_PT_FSM47  (KNN_DATA_PT_CORE47),


	.KNN_DATA_PT_FSM48  (KNN_DATA_PT_CORE48),
	.KNN_DATA_PT_FSM49  (KNN_DATA_PT_CORE49),
	.KNN_DATA_PT_FSM50  (KNN_DATA_PT_CORE50),
	.KNN_DATA_PT_FSM51  (KNN_DATA_PT_CORE51),
	.KNN_DATA_PT_FSM52  (KNN_DATA_PT_CORE52),
	.KNN_DATA_PT_FSM53  (KNN_DATA_PT_CORE53),
	.KNN_DATA_PT_FSM54  (KNN_DATA_PT_CORE54),
	.KNN_DATA_PT_FSM55  (KNN_DATA_PT_CORE55),
	
	.KNN_DATA_PT_FSM56  (KNN_DATA_PT_CORE56),
	.KNN_DATA_PT_FSM57  (KNN_DATA_PT_CORE57),
	.KNN_DATA_PT_FSM58  (KNN_DATA_PT_CORE58),
	.KNN_DATA_PT_FSM59  (KNN_DATA_PT_CORE59),
	.KNN_DATA_PT_FSM60  (KNN_DATA_PT_CORE60),
	.KNN_DATA_PT_FSM61  (KNN_DATA_PT_CORE61),
	.KNN_DATA_PT_FSM62  (KNN_DATA_PT_CORE62),
	.KNN_DATA_PT_FSM63  (KNN_DATA_PT_CORE63),
	
	.KNN_DATA_PT_FSM64  (KNN_DATA_PT_CORE64),
	.KNN_DATA_PT_FSM65  (KNN_DATA_PT_CORE65),
	.KNN_DATA_PT_FSM66  (KNN_DATA_PT_CORE66),
	.KNN_DATA_PT_FSM67  (KNN_DATA_PT_CORE67),
	.KNN_DATA_PT_FSM68  (KNN_DATA_PT_CORE68),
	.KNN_DATA_PT_FSM69  (KNN_DATA_PT_CORE69),
	.KNN_DATA_PT_FSM70  (KNN_DATA_PT_CORE70),
	.KNN_DATA_PT_FSM71  (KNN_DATA_PT_CORE71),
	
	.KNN_DATA_PT_FSM72  (KNN_DATA_PT_CORE72),
	.KNN_DATA_PT_FSM73  (KNN_DATA_PT_CORE73),
	.KNN_DATA_PT_FSM74  (KNN_DATA_PT_CORE74),
	.KNN_DATA_PT_FSM75  (KNN_DATA_PT_CORE75),
	.KNN_DATA_PT_FSM76  (KNN_DATA_PT_CORE76),
	.KNN_DATA_PT_FSM77  (KNN_DATA_PT_CORE77),
	.KNN_DATA_PT_FSM78  (KNN_DATA_PT_CORE78),
	.KNN_DATA_PT_FSM79  (KNN_DATA_PT_CORE79),
	
	.KNN_DATA_PT_FSM80  (KNN_DATA_PT_CORE80),
	.KNN_DATA_PT_FSM81  (KNN_DATA_PT_CORE81),
	.KNN_DATA_PT_FSM82  (KNN_DATA_PT_CORE82),
	.KNN_DATA_PT_FSM83  (KNN_DATA_PT_CORE83),
	.KNN_DATA_PT_FSM84  (KNN_DATA_PT_CORE84),
	.KNN_DATA_PT_FSM85  (KNN_DATA_PT_CORE85),
	.KNN_DATA_PT_FSM86  (KNN_DATA_PT_CORE86),
	.KNN_DATA_PT_FSM87  (KNN_DATA_PT_CORE87),
	
	.KNN_DATA_PT_FSM88  (KNN_DATA_PT_CORE88),
	.KNN_DATA_PT_FSM89  (KNN_DATA_PT_CORE89),
	.KNN_DATA_PT_FSM90  (KNN_DATA_PT_CORE90),
	.KNN_DATA_PT_FSM91  (KNN_DATA_PT_CORE91),
	.KNN_DATA_PT_FSM92  (KNN_DATA_PT_CORE92),
	.KNN_DATA_PT_FSM93  (KNN_DATA_PT_CORE93),
	.KNN_DATA_PT_FSM94  (KNN_DATA_PT_CORE94),
	.KNN_DATA_PT_FSM95  (KNN_DATA_PT_CORE95),
	
	
	.KNN_DATA_PT_FSM96  (KNN_DATA_PT_CORE96),
	.KNN_DATA_PT_FSM97  (KNN_DATA_PT_CORE97),
	.KNN_DATA_PT_FSM98  (KNN_DATA_PT_CORE98),
	.KNN_DATA_PT_FSM99  (KNN_DATA_PT_CORE99),
	.KNN_DATA_PT_FSM100  (KNN_DATA_PT_CORE100),
	.KNN_DATA_PT_FSM101  (KNN_DATA_PT_CORE101),
	.KNN_DATA_PT_FSM102  (KNN_DATA_PT_CORE102),
	.KNN_DATA_PT_FSM103  (KNN_DATA_PT_CORE103),
	
	
	.KNN_DATA_PT_FSM104  (KNN_DATA_PT_CORE104),
	.KNN_DATA_PT_FSM105  (KNN_DATA_PT_CORE105),
	.KNN_DATA_PT_FSM106  (KNN_DATA_PT_CORE106),
	.KNN_DATA_PT_FSM107  (KNN_DATA_PT_CORE107),
	.KNN_DATA_PT_FSM108  (KNN_DATA_PT_CORE108),
	.KNN_DATA_PT_FSM109  (KNN_DATA_PT_CORE109),
	.KNN_DATA_PT_FSM110  (KNN_DATA_PT_CORE110),
	.KNN_DATA_PT_FSM111  (KNN_DATA_PT_CORE111),
	
	
	.KNN_DATA_PT_FSM112  (KNN_DATA_PT_CORE112),
	.KNN_DATA_PT_FSM113  (KNN_DATA_PT_CORE113),
	.KNN_DATA_PT_FSM114  (KNN_DATA_PT_CORE114),
	.KNN_DATA_PT_FSM115  (KNN_DATA_PT_CORE115),
	.KNN_DATA_PT_FSM116  (KNN_DATA_PT_CORE116),
	.KNN_DATA_PT_FSM117  (KNN_DATA_PT_CORE117),
	.KNN_DATA_PT_FSM118  (KNN_DATA_PT_CORE118),
	.KNN_DATA_PT_FSM119  (KNN_DATA_PT_CORE119),
	
	.KNN_DATA_PT_FSM120  (KNN_DATA_PT_CORE120),
	.KNN_DATA_PT_FSM121  (KNN_DATA_PT_CORE121),
	.KNN_DATA_PT_FSM122  (KNN_DATA_PT_CORE122),
	.KNN_DATA_PT_FSM123  (KNN_DATA_PT_CORE123),
	.KNN_DATA_PT_FSM124  (KNN_DATA_PT_CORE124),
	.KNN_DATA_PT_FSM125  (KNN_DATA_PT_CORE125),
	.KNN_DATA_PT_FSM126  (KNN_DATA_PT_CORE126),
	.KNN_DATA_PT_FSM127  (KNN_DATA_PT_CORE127),
	
	.KNN_TEST_PT_FSM  (KNN_TEST_PT_CORE),
	.KNN_VALID_IN_FSM (KNN_VALID_CORE),
	.KNN_VALID_O      (KNN_VALID_OUT_CORE),
	.clk(CLK_CORE),
	.rst(RST_CORE)
	);


//////////////////////////////////////////////////////////////////////////
knn_datapath knn_datapath_inst
(
	//from fsm
	 .KNN_TEST_PT_DP(KNN_TST_CORE),
	 .KNN_DATA_PT_DP(KNN_DAT_CORE),
	 .KNN_START_DP(KNN_ST_CORE),
	
	//from sw reg
	 .KNN_SAMPLE_DP(KNN_SAMPLE_CORE),
	//to sw reg
	.KN1_OUT(KN1_OUT_CORE),
	.KN2_OUT(KN2_OUT_CORE),
	.KN3_OUT(KN3_OUT_CORE),
	.KN4_OUT(KN4_OUT_CORE),
	.KN5_OUT(KN5_OUT_CORE),
	.KN6_OUT(KN6_OUT_CORE),
	
	.IN1_OUT(IN1_OUT_CORE),
	.IN2_OUT(IN2_OUT_CORE),
	.IN3_OUT(IN3_OUT_CORE),
	.IN4_OUT(IN4_OUT_CORE),
	.IN5_OUT(IN5_OUT_CORE),
	.IN6_OUT(IN6_OUT_CORE),
		
	.clk(CLK_CORE),
	.rst(RST_CORE)
);
		
endmodule 
